LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.mux16to1_package.all;
USE work.mux2to1_package.all;

ENTITY mux_32to1 IS
GENERIC (N : INTEGER := 32);
	PORT (S           					: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			X0,X1,X2,X3,X4,X5,X6,X7,X8	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X9,X10,X11,X12,X13,X14,X15	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X16,X17,X18,X19,X20,X21,X22: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X23,X24,X25,X26,X27,X28,X29: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X30,X31							: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			Y									: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END mux_32to1;

ARCHITECTURE Structure OF mux_32to1 IS
	SIGNAL W0,W1	: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN
	MUX0_16_1:	mux_16to1 PORT MAP(S(0),S(1),S(2),S(3),X0,X1,X2,X3,X4,X5,X6,
												X7,X8,X9,X10,X11,X12,X13,X14,X15,W0);
												
	MUX1_16_1:	mux_16to1 PORT MAP(S(0),S(1),S(2),S(3),X16,X17,X18,X19,X20,X21,
											 X22,X23,X24,X25,X26,X27,X28,X29,X30,X31,W1);
											 
	MUX2_2_1	:	mux_2to1 GENERIC MAP(N) PORT MAP(S(4),W0,W1,Y);
END Structure;
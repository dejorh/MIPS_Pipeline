LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.mux8to1_package.all;
USE work.mux2to1_package.all;

ENTITY mux_16to1 IS
GENERIC (N : INTEGER := 32);
	PORT (S0,S1,S2,S3		: IN STD_LOGIC;
			X0,X1,X2,X3		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X4,X5,X6,X7		: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X8,X9,X10,X11	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			X12,X13,X14,X15: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			Y					: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END mux_16to1;

ARCHITECTURE Structure OF mux_16to1 IS
	SIGNAL W0,W1	: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN
	MUX0_8_1	:	mux_8to1	PORT MAP(S0,S1,S2,X0,X1,X2,X3,X4,X5,X6,X7,W0);
	MUX1_8_1	:	mux_8to1 PORT MAP(S0,S1,S2,X8,X9,X10,X11,X12,X13,X14,X15,W1);
	MUX2_2_1	:	mux_2to1 GENERIC MAP(N) PORT MAP(S3,W0,W1,Y);
END Structure;
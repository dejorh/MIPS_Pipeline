LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.mux2to1_package.all;

ENTITY mux_4to1 IS
GENERIC (N : INTEGER := 32);
	PORT (S				: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			X0,X1,X2,X3	: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			Y				: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END mux_4to1;

ARCHITECTURE Structure OF mux_4to1 IS
	SIGNAL W0,W1	: STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN
	MUX0_2_1	:	mux_2to1	GENERIC MAP(N) PORT MAP(S(0),X0,X1,W0);
	MUX1_2_1	:	mux_2to1 GENERIC MAP(N) PORT MAP(S(0),X2,X3,W1);
	MUX2_2_1	:	mux_2to1 GENERIC MAP(N) PORT MAP(S(1),W0,W1,Y);
END Structure;
LIBRARY ieee;						--Provide compiler with access to Library
USE ieee.std_logic_1164.all;	--Use all contents from package in ieee Library

PACKAGE HDU_1_package IS
	COMPONENT Hazard_Detect					--Component Declaration
	GENERIC(M : INTEGER := 5);
		PORT (EX_MEM_PCSrc: IN STD_LOGIC;
				ID_EX_MemRead,ID_EX_Jump	: IN STD_LOGIC;
				IF_ID_Rs,IF_ID_Rt,ID_EX_Rt	: IN STD_LOGIC_VECTOR(M-1 DOWNTO 0);
				PC_Write,IF_ID_Write,Flush	: OUT STD_LOGIC);
	END COMPONENT;
END HDU_1_package;
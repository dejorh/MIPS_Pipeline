LIBRARY ieee;							--Provide compiler with access to Library
USE ieee.std_logic_1164.all;		--Use all contents from package in ieee Library

PACKAGE Reg32en_package IS
	COMPONENT Reg32en						--Component Declaration
		GENERIC(N	: INTEGER := 32);	-- Constant declaration
		PORT (En,Clock,Reset	:  IN  STD_LOGIC;				--Input declaration
			D					:	IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				--Output declaration
			Q					:	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
	END COMPONENT;
END Reg32en_package;
LIBRARY ieee;						--Provide compiler with access to Library
USE ieee.std_logic_1164.all;	--Use all contents from package in ieee Library

PACKAGE IExecute_package IS
	COMPONENT IExecute_Stage			--Component Declaration
		GENERIC(N  : INTEGER := 32);	-- Constant declaration
					--select read_data_2 for R-Type and Sign-Extend value for I-Type
		PORT (ALU_Src						: IN STD_LOGIC; 
					-- Select Vector for ALU operations
				ALU_ctrl						: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
						-- Data to be read from read registers
				read_data_1					: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
				read_data_2					: BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0);
						-- The Sign-Extended value
				Extend_value				: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
						-- ALU output
				ALU_result					: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
						-- Zero signal, also an ouput
				Zero							: OUT STD_LOGIC);
	END COMPONENT;
END IExecute_package;